`ifndef __rename_intf
`define __rename_intf

interface rename_interface_dut;
  logic        clk;
  logic        valid; 
  logic  [2:0] addr;
  logic        irq; 

 import uvm_pkg::*;
      
//ASERTII
      
endinterface


`endif